package axi_test_pkg;

        import uvm_pkg::*;

        `include "uvm_macros.svh"
        `include "axi_xtn.sv"
        `include "axi_m_agt_config.sv"
        `include "axi_s_agt_config.sv"
        `include "axi_env_config.sv"
        `include "axi_m_drv.sv"
        `include "axi_m_mon.sv"
        `include "axi_m_seqr.sv"
        `include "axi_m_agt.sv"
        `include "axi_m_agt_top.sv"
        `include "axi_m_seq.sv"
        `include "axi_s_drv.sv"
        `include "axi_s_mon.sv"
        `include "axi_s_seqr.sv"
        `include "axi_s_agt.sv"
        `include "axi_s_agt_top.sv"
        `include "axi_s_seq.sv"
        `include "axi_v_seqr.sv"
        `include "axi_v_seqs.sv"
        `include "axi_sb.sv"
        `include "axi_interconnect.sv"
        `include "axi_env.sv"
        //`include "axi_interconnect.sv"
        `include "axi_base_test.sv"
        //`include "axi_interconnect.sv"

endpackage

